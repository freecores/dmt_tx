

`define VENDOR_FPGA


